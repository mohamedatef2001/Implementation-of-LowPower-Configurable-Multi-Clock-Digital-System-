module BIT_SYNC_TB #(parameter NUM_STG_TB = 3 ,DEPTH_TB   = 3 )();
reg                           CLK_TB      ;
reg                           RST_TB     ;
reg      [DEPTH_TB-1:0]       ASYNC_TB   ;
wire     [DEPTH_TB-1:0]       SYNC_TB    ;

  
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 ////////////  PARAMETERS ///////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/

parameter CLK_P     = 10 ;
                    
          
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 //////////// INSTANTIATION /////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                 
					 
BIT_SYNC  # ( .NUM_STG(NUM_STG_TB) , .DEPTH(DEPTH_TB) )  DUT
(
.clk(CLK_TB),
.rst(RST_TB),
.async(ASYNC_TB),
.sync(SYNC_TB)
);

                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 /////////////// CLOCK //////////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                 
               
 always  #(CLK_P/2) CLK_TB = ~ CLK_TB; 
 
 
 
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 //////////// INITIAL BLOCK /////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                             
initial
begin
      $dumpfile("UART_RX_TB.vcd");
      $dumpvars;
      initialize();
      ASYNC_TB = 'b101;
     #25
     ASYNC_TB = 'b010;
     #100
     $finish;  // CHECK WAVEFORM
end
      
 
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 //////////////// TASKS /////////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                 
      
 task initialize ;                                      // IDEAL STATE
  begin
        //#(CLK_P);
        CLK_TB = 'b0;
        RST_TB = 'b0;
        #(CLK_P);
        RST_TB = 'b1;
        //#(CLK_P);
  end
endtask     


endmodule

