module RST_SYNC_TB #(parameter NUM_STG_TB = 3) ();
reg                 CLK_TB ;
reg                 RST_TB ;
wire                SYNC_RST_TB ;



  
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 ////////////  PARAMETERS ///////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/

parameter CLK_P     = 10 ;
                    
          
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 //////////// INSTANTIATION /////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                 
					 
RST_SYNC  # ( .NUM_STG(NUM_STG_TB) )  DUT
(
.clk(CLK_TB),
.rst(RST_TB),
.sync_rst(SYNC_RST_TB)
);

                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 /////////////// CLOCK //////////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                 
               
 always  #(CLK_P/2) CLK_TB = ~ CLK_TB; 
 
 
 
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 //////////// INITIAL BLOCK /////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                             
initial
begin
      $dumpfile("UART_RX_TB.vcd");
      $dumpvars;
      initialize();
      RST_TB = 'b0;
      #8
      RST_TB = 'b1;
      #100
     $finish;  // CHECK WAVEFORM
end
      
 
                 /*//////////////////////////////////////
                 ////////////////////////////////////////
                 //////////////// TASKS /////////////////
                 ////////////////////////////////////////
                 //////////////////////////////////////*/
                 
      
 task initialize ;                                      // IDEAL STATE
  begin
        CLK_TB = 'b0;
        RST_TB = 'b1;
        #(CLK_P);
        //RST_TB = 'b1;
  end
endtask     


endmodule



